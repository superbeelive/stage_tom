Inverse RIAA test circuit
v1 1 0 AC 1.0

r1 1 2 27k
r2 1 2 27k
c1 1 2 5.6n
r4 2 3 150k
c2 2 3 22n
r5 3 0 470

.ac dec 100 20 20000
.plot ac vdb(3)

* Commands for Spice3
*#run
*#plot db(v(3))
.end

