* PSpice current controlled switch example

C1 1 0 40UF IC=200
VX 2 1 DC 0V
W1 2 3 VX SMOD

.MODEL SMOD ISWITCH(RON=1E6 ROFF=0.001 ION=1MA IOFF=0)

L1 3 0 50UH

.TRAN 1US 160US UIC

.PLOT TRAN V(1) I(VX)
.PROBE
.END
