SIMPLE DIFFERENTIAL PAIR
.OPTIONS NOPAGE ACCT
.WIDTH OUT=80
.TEMP 50
.TRAN 2N 100N 
.PLOT  TRAN V(4) V(1)

VIN 1 0 PWL (0NS -.2V 10NS -.2V 14NS .2V 100NS .2V)
VCC 7 0  12
VEE 8 0 -12
*
Q1 3 2 4 QNL
Q2 5 6 4 QNL
*
RS1   1 2 1K
RS2   6 0 1K
RC1   3 7 10K
RC2   5 7 10K 
RBIAS 4 8 10K
*
.MODEL QNL NPN(BF=100 RB=100 CCS=2PF TF=0.3NS TR=6NS CJE=3PF CJC=2PF
+   VA=50)
.END
