Example 9.1 Output characteristics of N-channel JFET

.OPTION LIMPTS=500

* Gate to source voltage of 0V

VGS 1 0 DC 0V

* A dummy voltage source of 0V

VX 3 2 DC 0V

* DC supply voltage of 12V

VDD 3 0 DC 12V

* J1 with model JMOD

J1 2 1 0 JMOD

.MODEL JMOD NJF (IS=100e-14 RD=10 RS=10 BETA=1E-3 VTO=-5)

* VDD is swept from 0 to 12V and VGS from 0 to -4V.

.DC VDD 0 12 0.2 VGS 0 -4 1
.PLOT DC I(VX)

* Commands for Spice3
*#run
*#plot vx#branch

.END
