voltage divider netlist
V1 a 0 1
R1 a b 1k
R2 b 0 2k
.end
