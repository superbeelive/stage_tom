FM de-emphasis circuit (50us)
v1 1 0 AC 1.0
r1 1 2 5k
c1 2 0 10n
.ac dec 100 20 20000
.plot ac vdb(2)

* Commands for Spice3
*#run
*#plot v(2)
.end

