.exercice 2 
Vin in 0 dc 0 ac 1 sin(0 1m 50)
l1 in out 3
R1 out 0 1k
.end
