Example 10.7 Differential Amplifier

.WIDTH OUT=80

VCC  11  0  12V
VEE  0   10 12V
VIN  1   0  DC 0.25

RC1 11   3  10K
RC2 11   5  10K
RE1  4  12  150
RE2  7  12  150
RS1  1   2  1.5K
RS2  6   0  1.5K
RX  11   8  20K

Q1   3   2   4  QN
Q2   5   6   7  QN
Q3  12   8   9  QN
Q4   9   9  10  QN
Q5   8   9  10  QN


* DC transfer function analysis

.TF V(3,5) VIN


* Model for NPN BJTs with model name QN

.MODEL QN NPN (BF=50 RB=70 RC=40)
.END
